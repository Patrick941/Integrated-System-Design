module scoreboard(
    input clk,
    input reset
);

    initial begin
        $display("scoreboard: Starting simulation");
    end


endmodule